module gate(
input a,
input b,

output z
);

or (z, a, b);

endmodule