module try;
initial
begin
	$display ("This is a simple code");
	$finish;
end
endmodule