module GreenRoad;
  initial 
    begin
      $display("Learning Verilog is easy");
      $finish ;
    end
endmodule